//Gate Level
module mynotgate(
    input wire a,
    output wire nota
);


not inv1(nota,a); // Inverter gate

endmodule