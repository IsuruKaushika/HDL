module myfirstprog ();

    initial begin
        $display("Hello");
        $finish;
    end
endmodule