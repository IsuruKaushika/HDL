module mynotgate(
    input wire a,
    output wire nota
    );

assign nota =~a;

endmodule

//RTL